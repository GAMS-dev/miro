header 1|header 2|Value 1|header 4|Value 2
j1|i1|12.34|bla1|1
j2|i2|13.470|bla2|2
j3|i3|16.471|bla3|3
j4|i4|11|bla4|4
j5|i5|13.477|bla5|5
j6|i6|7|bla6|6
j7|i7|13.4791|bla7|7
